`include "uvm.sv"
`include "uvm_macros.svh"
import  uvm_pkg::*;

`include "WB2APB_interface.sv"
`include "WB2APB_seq_item.sv"
`include "WB2APB_sequence.sv"
`include "WB2APB_sequencer.sv"
`include "WB2APB_driver.sv"
`include "WB2APB_monitor.sv"
`include "WB2APB_agent.sv"
`include "WB2APB_scoreboard.sv"
`include "WB2APB_env.sv"
`include "WB2APB_sva.sv"


`include "WB2APB_base_test.sv"
`include "WB2APB_test.sv"